entity CMDBUFFERS is 
port(

);
end CMDBUFFERS

architecture CMDBUFFERS_Arch of CMDBUFFERS is
begin
    